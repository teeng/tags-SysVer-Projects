/*
Constructs a 16x1 multiplexer module named mux16_1
	out is the output for the mux with type logic
	in is 16'b input for the mux with type logic
	sel is 4'b select line for the mux with type logic
	
	Timescale was a necessary addition to the module for running
		given regstim simulation file without errors.
*/
`timescale 1 ps / 1 ps

module mux16_1(out, in, sel);
	output logic out;
	input  logic [15:0] in;
	input logic [3:0] sel;
	
	// internal logic 2'b v is to store
		// results of two of the two 8x1 muxes needed to determine the final
		// 16x1 mux output
	logic  [1:0] v;
	// instantiates two 8x1 mux8_1 named m2, m1.
	// m2 and m1 both have outputs to the internal signals v0 and v1,1
		// where the 2'b combined result is used in a 3rd mux2_1, m0.
	// m2 and m1 are controlled by the 0th to 2nd bit from the select line, sel
	// m0 uses the 3rd bit from the select line, sel, with output out for the mux16_1 module.
	mux8_1 m2 (.out(v[0]),  .in(in[7:0]), .sel(sel[2:0]));
	mux8_1 m1 (.out(v[1]),  .in(in[15:8]), .sel(sel[2:0])); 
	mux2_1 m0 (.out(out), .in(v),  .sel(sel[3]));
endmodule

module mux16_1_testbench();
	logic [15:0] in;
	logic [3:0] sel;    
	logic  out;
	
	mux16_1 dut (.out, .in, .sel);
	
	integer i;   
	initial begin  
		for(i=0; i<8; i++) begin  
			{sel, in} = i; #3000;
		end
		
		sel <= 4'b0001;
		for(i=0; i<8; i++) begin  
			in = i; #3000;
		end
		
		sel <= 4'b0010;
		for(i=0; i<8; i++) begin  
			in = i; #3000;
		end
		
		sel <= 4'b0011;
		for(i=0; i<16; i++) begin  
			in = i; #3000;
		end
		
	$stop;
	end  
endmodule 